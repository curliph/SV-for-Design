module asymmetric_ram #(
) (
);

endmodule
