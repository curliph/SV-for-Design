// ADD/SUB Design {SUB = using 2's Complement Addition}
module optimal_add_sub #(
) (
);

endmodule
