module interrupt_controller #(
) (
  input  logic clk,
  input  logic reset,
);

endmodule
