module jtag_tap_controller #(
) (
);

endmodule
