module cpu_mx1_interconnect #(
) (
);

endmodule
