module data_mux #(
) (
);

endmodule

module data_demux #(
) (
);

endmodule
