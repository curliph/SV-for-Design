module freq_comparator #(
  parameter DATA_WIDTH = 32
) (
);

endmodule
